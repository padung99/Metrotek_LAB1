module top_tb;

bit_population_counter_tb #(.WIDTH_TB(5)) dut1 ();
bit_population_counter_tb #(.WIDTH_TB(10)) dut2 ();
bit_population_counter_tb #(.WIDTH_TB(16)) dut3 ();

endmodule